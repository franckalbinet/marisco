netcdf maris {
// Custom types
types:
  int64 enum area_t {TBD_1 = 0} ;
  int64 enum bio_group_t {TBD_2 = 0} ;
  int64 enum body_part_t {TBD_3 = 0} ;
  int64 enum count_met_t {TBD_4 = 0} ;
  int64 enum dl_t {TBD_5 = 0} ;
  int64 enum filt_t {TBD_6 = 0} ;
  int64 enum nuclide_t {TBD_7 = 0} ;
  int64 enum prep_met_t {TBD_8 = 0} ;
  int64 enum samp_met_t {TBD_9 = 0} ;
  int64 enum sed_type_t {TBD_10 = 0} ;
  int64 enum species_t {TBD_11 = 0} ;
  int64 enum unit_t {TBD_12 = 0} ;
  int64 enum lab_t {TBD_13 = 0};
    
// Global attributes
:id = "TBD" ;
:title = "TBD" ;
:summary = "TBD" ;  
:keywords = "TBD" ;
:history = "TBD" ; // ex: "Created 2024" ;
:keywords_vocabulary = "GCMD Science Keywords" ;
:keywords_vocabulary_url = "https://gcmd.earthdata.nasa.gov/static/kms/" ;
:record = "TBD" ;
:featureType = "TBD" ;
:cdm_data_type = "TBD" ;
:Conventions = "CF-1.10 ACDD-1.3" ;
:publisher_name = "Paul MCGINNITY, Iolanda OSVATH, Florence DESCROIX-COMANDUCCI" ;
:publisher_email = "p.mc-ginnity@iaea.org, i.osvath@iaea.org, F.Descroix-Comanducci@iaea.org" ;
:publisher_url = "https://maris.iaea.org" ;
:publisher_institution = "International Atomic Energy Agency - IAEA" ;
:creator_name = "TBD" ;
:institution = "TBD" ;
:metadata_link = "TBD" ;
:creator_email = "TBD" ;
:creator_url = "TBD" ;
:references = "TBD" ;
:license = "Without prejudice to the applicable Terms and Conditions (https://nucleus.iaea.org/Pages/Others/Disclaimer.aspx), I hereby agree that any use of the data will contain appropriate acknowledgement of the data source(s) and the IAEA Marine Radioactivity Information System (MARIS)." ;
:comment = "TBD" ;
:geospatial_lat_min = "TBD" ;
:geospatial_lon_min = "TBD" ;
:geospatial_lat_max = "TBD" ;
:geospatial_lon_max = "TBD" ;
:geospatial_vertical_min = "TBD" ;
:geospatial_vertical_max = "TBD" ;
:geospatial_bounds = "TBD" ;
:geospatial_bounds_crs = "EPSG:4326" ;
:time_coverage_start = "TBD" ;
:time_coverage_end = "TBD" ;
:local_time_zone = "TBD" ;
:date_created = "TBD" ;
:date_modified = "TBD" ;
:publisher_postprocess_logs = "TBD" ; // Logs of the processing steps

// Root dimension
//dimensions:
//    id = UNLIMITED ;

// Groups
group: biota {  
    dimensions:
        id = UNLIMITED ;
    variables:
        // Common variables
        uint64 id(id) ;
            id:long_name = "Measurement ID" ;
        float lon(id) ;   
            lon:long_name = "Measurement longitude" ;
            lon:standard_name = "longitude" ;
            lon:units = "degrees_east" ;
        float lat(id) ;
            lat:long_name = "Measurement latitude" ;
            lat:standard_name = "latitude" ;
            lat:units = "degrees_north" ;
        float smp_depth(id) ;
            smp_depth:long_name = "Sample depth below seal level" ;
            smp_depth:standard_name = "sample_depth_below_sea_floor" ;
            smp_depth:units = "m" ;
            smp_depth:axis = "Z" ;
        float tot_depth(id) ;
            tot_depth:long_name = "Total depth below seal level" ;
            tot_depth:standard_name = "total_depth_below_sea_floor" ;
            tot_depth:units = "m" ;
            tot_depth:axis = "Z" ;
        uint64 time(id) ;
            time:long_name = "Time of measurement" ;
            time:standard_name = "time" ;
            time:units = "seconds since 1970-01-01 00:00:00.0" ;
            time:time_origin = "1970-01-01 00:00:00" ;
            time:time_zone = "UTC" ;
            time:abbreviation = "Date/Time" ;
            time:axis = "T" ;
            time:calendar = "gregorian" ;
        area_t area(id) ;
            area:long_name = "Marine area/region id" ;
            area:standard_name = "area_id" ;
        uint64 smp_id(id) ;
            smp_id:long_name = "Data provider sample ID" ;
            smp_id:standard_name = "sample_id" ;
        nuclide_t nuclide(id) ;
            nuclide:long_name = "Nuclide" ;
            nuclide:standard_name = "nuclide" ;
        float value(id) ;
            value:long_name = "Activity" ;
            value:standard_name = "activity" ;
        unit_t unit(id) ;
            unit:long_name = "Unit" ;
            unit:standard_name = "unit" ;
        float unc(id) ;
            unc:long_name = "Uncertainty" ;
            unc:standard_name = "uncertainty" ;
        dl_t dl(id) ;
            dl:long_name = "Detection limit" ;
            dl:standard_name = "detection_limit" ;
        filt_t filt(id) ;
            filt:long_name = "Filtering method" ;
            filt:standard_name = "filtered" ;
        count_met_t count_met(id) ;
            count_met:long_name = "Counting method" ;
            count_met:standard_name = "counting_method" ;
        samp_met_t samp_met(id) ;
            samp_met:long_name = "Sampling method" ;
            samp_met:standard_name = "sampling_method" ;
        prep_met_t prep_met(id) ;
            prep_met:long_name = "Preparation method" ;
            prep_met:standard_name = "preparation_method" ;
        lab_t lab(id) ;
            lab:long_name = "laboratory" ;
            lab:standard_name = "laboratory" ;
        float vol(id) ;
            vol:long_name = "Volume" ;
            vol:standard_name = "volume" ;
        float sal(id) ;
            sal:long_name = "Salinity" ;
            sal:standard_name = "salinity" ;
        float temp(id) ;
            temp:long_name = "Temperature" ;
            temp:standard_name = "temperature" ;
        float ph(id) ;
            ph:long_name = "pH" ;
            ph:standard_name = "pH" ;

        // Biota specific variables
        bio_group_t bio_group(id) ;
            bio_group:long_name = "Biota group" ;
            bio_group:standard_name = "biota_group_tbd" ;
        species_t species(id) ;
            species:long_name = "Species" ;
            species:standard_name = "species" ;
        body_part_t body_part(id) ;
            body_part:long_name = "Body part" ;
            body_part:standard_name = "body_part_tbd" ;
		float drywt(id) ;
        	drywt:long_name = "Dry weight of biota sample, expressed in grams." ;
        	drywt:standard_name = "dry_weight_of_biota_sample" ;
		float wetwt(id) ;
            wetwt:long_name = "Wet weight of biota sample, expressed in grams." ;
            wetwt:standard_name = "wet_weight_of_biota_sample" ;
		float percentwt(id) ;
        	percentwt:long_name = "Dry weight as a percentage of fresh weight." ;
        	percentwt:standard_name = "percentage_weight_of_biota_sample" ;
}

group: seawater {
    dimensions:
        id = UNLIMITED ;
    variables:
        // Common variables
        uint64 id(id) ;
            id:long_name = "Measurement ID" ;
        float lon(id) ;   
            lon:long_name = "Measurement longitude" ;
            lon:standard_name = "longitude" ;
            lon:units = "degrees_east" ;
        float lat(id) ;
            lat:long_name = "Measurement latitude" ;
            lat:standard_name = "latitude" ;
            lat:units = "degrees_north" ;
        float smp_depth(id) ;
            smp_depth:long_name = "Sample depth below seal level" ;
            smp_depth:standard_name = "sample_depth_below_sea_floor" ;
            smp_depth:units = "m" ;
            smp_depth:axis = "Z" ;
        float tot_depth(id) ;
            tot_depth:long_name = "Total depth below seal level" ;
            tot_depth:standard_name = "total_depth_below_sea_floor" ;
            tot_depth:units = "m" ;
            tot_depth:axis = "Z" ;
        uint64 time(id) ;
            time:long_name = "Time of measurement" ;
            time:standard_name = "time" ;
            time:units = "seconds since 1970-01-01 00:00:00.0" ;
            time:time_origin = "1970-01-01 00:00:00" ;
            time:time_zone = "UTC" ;
            time:abbreviation = "Date/Time" ;
            time:axis = "T" ;
            time:calendar = "gregorian" ;
        area_t area(id) ;
            area:long_name = "Marine area/region id" ;
            area:standard_name = "area_id" ;
        uint64 smp_id(id) ;
            smp_id:long_name = "Data provider sample ID" ;
            smp_id:standard_name = "sample_id" ;
        nuclide_t nuclide(id) ;
            nuclide:long_name = "Nuclide" ;
            nuclide:standard_name = "nuclide" ;
        float value(id) ;
            value:long_name = "Activity" ;
            value:standard_name = "activity" ;
        unit_t unit(id) ;
            unit:long_name = "Unit" ;
            unit:standard_name = "unit" ;
        float unc(id) ;
            unc:long_name = "Uncertainty" ;
            unc:standard_name = "uncertainty" ;
        dl_t dl(id) ;
            dl:long_name = "Detection limit" ;
            dl:standard_name = "detection_limit" ;
        filt_t filt(id) ;
            filt:long_name = "Filtering method" ;
            filt:standard_name = "filtered" ;
        count_met_t count_met(id) ;
            count_met:long_name = "Counting method" ;
            count_met:standard_name = "counting_method" ;
        samp_met_t samp_met(id) ;
            samp_met:long_name = "Sampling method" ;
            samp_met:standard_name = "sampling_method" ;
        prep_met_t prep_met(id) ;
            prep_met:long_name = "Preparation method" ;
            prep_met:standard_name = "preparation_method" ;
        lab_t lab(id) ;
            lab:long_name = "laboratory" ;
            lab:standard_name = "laboratory" ;
        float vol(id) ;
            vol:long_name = "Volume" ;
            vol:standard_name = "volume" ;
        float sal(id) ;
            sal:long_name = "Salinity" ;
            sal:standard_name = "salinity" ;
        float temp(id) ;
            temp:long_name = "Temperature" ;
            temp:standard_name = "temperature" ;
        float ph(id) ;
            ph:long_name = "pH" ;
            ph:standard_name = "pH" ;
}

group: sediment {
    dimensions:
        id = UNLIMITED ;
    variables:
        // Common variables
        uint64 id(id) ;
            id:long_name = "Measurement ID" ;
        float lon(id) ;   
            lon:long_name = "Measurement longitude" ;
            lon:standard_name = "longitude" ;
            lon:units = "degrees_east" ;
        float lat(id) ;
            lat:long_name = "Measurement latitude" ;
            lat:standard_name = "latitude" ;
            lat:units = "degrees_north" ;
        float smp_depth(id) ;
            smp_depth:long_name = "Sample depth below seal level" ;
            smp_depth:standard_name = "sample_depth_below_sea_floor" ;
            smp_depth:units = "m" ;
            smp_depth:axis = "Z" ;
        float tot_depth(id) ;
            tot_depth:long_name = "Total depth below seal level" ;
            tot_depth:standard_name = "total_depth_below_sea_floor" ;
            tot_depth:units = "m" ;
            tot_depth:axis = "Z" ;
        uint64 time(id) ;
            time:long_name = "Time of measurement" ;
            time:standard_name = "time" ;
            time:units = "seconds since 1970-01-01 00:00:00.0" ;
            time:time_origin = "1970-01-01 00:00:00" ;
            time:time_zone = "UTC" ;
            time:abbreviation = "Date/Time" ;
            time:axis = "T" ;
            time:calendar = "gregorian" ;
        area_t area(id) ;
            area:long_name = "Marine area/region id" ;
            area:standard_name = "area_id" ;
        uint64 smp_id(id) ;
            smp_id:long_name = "Data provider sample ID" ;
            smp_id:standard_name = "sample_id" ;
        nuclide_t nuclide(id) ;
            nuclide:long_name = "Nuclide" ;
            nuclide:standard_name = "nuclide" ;
        float value(id) ;
            value:long_name = "Activity" ;
            value:standard_name = "activity" ;
        unit_t unit(id) ;
            unit:long_name = "Unit" ;
            unit:standard_name = "unit" ;
        float unc(id) ;
            unc:long_name = "Uncertainty" ;
            unc:standard_name = "uncertainty" ;
        dl_t dl(id) ;
            dl:long_name = "Detection limit" ;
            dl:standard_name = "detection_limit" ;
        filt_t filt(id) ;
            filt:long_name = "Filtering method" ;
            filt:standard_name = "filtered" ;
        count_met_t count_met(id) ;
            count_met:long_name = "Counting method" ;
            count_met:standard_name = "counting_method" ;
        samp_met_t samp_met(id) ;
            samp_met:long_name = "Sampling method" ;
            samp_met:standard_name = "sampling_method" ;
        prep_met_t prep_met(id) ;
            prep_met:long_name = "Preparation method" ;
            prep_met:standard_name = "preparation_method" ;
        lab_t lab(id) ;
            lab:long_name = "laboratory" ;
            lab:standard_name = "laboratory" ;
        float vol(id) ;
            vol:long_name = "Volume" ;
            vol:standard_name = "volume" ;
        float sal(id) ;
            sal:long_name = "Salinity" ;
            sal:standard_name = "salinity" ;
        float temp(id) ;
            temp:long_name = "Temperature" ;
            temp:standard_name = "temperature" ;
        float ph(id) ;
            ph:long_name = "pH" ;
            ph:standard_name = "pH" ;

        // Sediment specific variables
        sed_type_t sed_type(id) ;
            sed_type:long_name = "Sediment type" ;
            sed_type:standard_name = "sediment_type_tbd" ;  
        float top(id) ;
            top:long_name = "Top depth of sediment layer" ;
            top:standard_name = "top_depth_of_sediment_layer_tbd" ;
        float bottom(id) ;
            bottom:long_name = "Bottom depth of sediment layer" ;
            bottom:standard_name = "bottom_depth_of_sediment_layer_tbd" ;
		float drywt(id) ;
            drywt:long_name = "Dry weight of sediment sample, expressed in grams." ;
            drywt:standard_name = "dry_weight_of_sediment_sample" ;
		float wetwt(id) ;
            wetwt:long_name = "Wet weight of sediment sample, expressed in grams." ;
            wetwt:standard_name = "wet_weight_of_sediment_sample" ;
		float percentwt(id) ;
        	percentwt:long_name = "Dry weight as a percentage of fresh weight." ;
        	percentwt:standard_name = "percentage_weight_of_biota_sample" ;
}

group: suspended_matter {
    dimensions:
        id = UNLIMITED ;
    variables:
        uint64 id(id) ;
            id:long_name = "Measurement ID" ;
        float lon(id) ;   
            lon:long_name = "Measurement longitude" ;
            lon:standard_name = "longitude" ;
            lon:units = "degrees_east" ;
        float lat(id) ;
            lat:long_name = "Measurement latitude" ;
            lat:standard_name = "latitude" ;
            lat:units = "degrees_north" ;
        float smp_depth(id) ;
            smp_depth:long_name = "Sample depth below seal level" ;
            smp_depth:standard_name = "sample_depth_below_sea_floor" ;
            smp_depth:units = "m" ;
            smp_depth:axis = "Z" ;
        float tot_depth(id) ;
            tot_depth:long_name = "Total depth below seal level" ;
            tot_depth:standard_name = "total_depth_below_sea_floor" ;
            tot_depth:units = "m" ;
            tot_depth:axis = "Z" ;
        uint64 time(id) ;
            time:long_name = "Time of measurement" ;
            time:standard_name = "time" ;
            time:units = "seconds since 1970-01-01 00:00:00.0" ;
            time:time_origin = "1970-01-01 00:00:00" ;
            time:time_zone = "UTC" ;
            time:abbreviation = "Date/Time" ;
            time:axis = "T" ;
            time:calendar = "gregorian" ;
        area_t area(id) ;
            area:long_name = "Marine area/region id" ;
            area:standard_name = "area_id" ;
        uint64 smp_id(id) ;
            smp_id:long_name = "Data provider sample ID" ;
            smp_id:standard_name = "sample_id" ;
        nuclide_t nuclide(id) ;
            nuclide:long_name = "Nuclide" ;
            nuclide:standard_name = "nuclide" ;
        float value(id) ;
            value:long_name = "Activity" ;
            value:standard_name = "activity" ;
        unit_t unit(id) ;
            unit:long_name = "Unit" ;
            unit:standard_name = "unit" ;
        float unc(id) ;
            unc:long_name = "Uncertainty" ;
            unc:standard_name = "uncertainty" ;
        dl_t dl(id) ;
            dl:long_name = "Detection limit" ;
            dl:standard_name = "detection_limit" ;
        filt_t filt(id) ;
            filt:long_name = "Filtering method" ;
            filt:standard_name = "filtered" ;
        count_met_t count_met(id) ;
            count_met:long_name = "Counting method" ;
            count_met:standard_name = "counting_method" ;
        samp_met_t samp_met(id) ;
            samp_met:long_name = "Sampling method" ;
            samp_met:standard_name = "sampling_method" ;
        prep_met_t prep_met(id) ;
            prep_met:long_name = "Preparation method" ;
            prep_met:standard_name = "preparation_method" ;
        lab_t lab(id) ;
            lab:long_name = "laboratory" ;
            lab:standard_name = "laboratory" ;
        float vol(id) ;
            vol:long_name = "Volume" ;
            vol:standard_name = "volume" ;
        float sal(id) ;
            sal:long_name = "Salinity" ;
            sal:standard_name = "salinity" ;
        float temp(id) ;
            temp:long_name = "Temperature" ;
            temp:standard_name = "temperature" ;
        float ph(id) ;
            ph:long_name = "pH" ;
            ph:standard_name = "pH" ;
}
}

netcdf enums_example {
    types:
        byte enum cloud_t {Clear = 0, Cumulonimbus = 1, Stratus = 2, 
            Stratocumulus = 3, Cumulus = 4, Altostratus = 5, Nimbostratus = 6, 
            Altocumulus = 7, Cirrostratus = 8, Cirrocumulus = 9, Cirrus = 10, 
            Missing = 127} ;

        byte enum sea_t {Clear = 0, Cumulonimbus = 1, Stratus = 2, 
            Stratocumulus = 3, Cumulus = 4, Altostratus = 5, Nimbostratus = 6, 
            Altocumulus = 7, Cirrostratus = 8, Cirrocumulus = 9, Cirrus = 10, 
            Missing = 127} ;

dimensions:
	time = UNLIMITED ; // (5 currently)
variables:
	cloud_t primary_cloud(time) ;
	    cloud_t primary_cloud:_FillValue = Missing ;

    sea_t primary_sea(time) ;
	    sea_t primary_sea:_FillValue = Missing ;
data:

 primary_cloud = Clear, Stratus, Clear, Cumulonimbus, _ ;
 primary_sea = Clear, Stratus, Clear, Cumulonimbus, _ ;
}